module portOR(
    input a, b, c,
    output d,
);

assign d = a & b & c;
endmodule
